library ieee;
use ieee.std_logic_1164.all;

library osvvm_common;
context osvvm_common.OsvvmCommonContext;
package AvalonStreamSlavePkg is
end package AvalonStreamSlavePkg;